
//
// module: p_mul_ftb
//
//  Dummy module for future use
//
module p_mul_ftb (
    input clock
    input resetn
);

endmodule
