
// TODO

module xc_sha256_ftb (

input clock,
input reset

);


endmodule
